`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Group:21
// Members: Debanjan Saha [19CS30014], Pritkumar Godhani [19CS10048]
//  
// Module Name: ShiftRegLeft 
// Project Name: Assignment-5 Question 4
//
//////////////////////////////////////////////////////////////////////////////////
module ShiftRegLeft(out, temp, data_in, clk, rst, load);
	input clk, load, rst;
	input [31:0] data_in;
	output reg out;
	output reg [31:0] temp;
	
	// Left Shift Logic + Asynchronous Load
	always @ (posedge clk or posedge load) begin
		if(load) 
			temp <= data_in;
		else if(rst)
			temp <= 16'b0;
		else begin
			out <= temp[31];
			temp <= {temp[30:0], 1'b0};
		end 
	end

endmodule 