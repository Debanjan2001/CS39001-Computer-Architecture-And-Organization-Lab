`include "rca64.v"

module TestRCA64();
    reg [63:0] a,b;
    reg cin;
    wire[63:0] sum;
    wire cout;

    RippleCarryAdder64 rca64(.A(a), .B(b), .cin(cin), .sum(sum), .cout(cout));

    initial begin
        $monitor("a = %b, b = %b, cin = %b, sum = %b, cout = %b", a, b, cin, sum, cout);
        #1 a = 64'b0000000000000000000000000000000011111111111111111111111111111111; b = 64'b0000000000000000000000000000000000000000000000000000000000000001; cin = 1'b0;
        #2 a = 64'b1111111111111111111111111111111111111111111111111111111111111111; b = 64'b0000000000000000000000000000000000000000000000000000000000000001; cin = 1'b0;
        #3 a = 64'b1111111111111111111111111111111111111111111111111111111111111111; b = 64'b0000000000000000000000000000000000000000000000000000000000000000; cin = 1'b1;
        #4 a = 64'b0000000000000001000000000000000100000000000000010000000000000001; b = 64'b0000000000000001000000000000000100000000000000010000000000000001; cin = 1'b0;
        #5 a = 64'b0010010011100001110001111100111101001000111000110101011000100111; b = 64'b0110101000111111100100100100111111111000100111110011111000100000; cin = 1'b0;
    end
endmodule